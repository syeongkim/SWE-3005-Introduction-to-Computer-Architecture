module testbench;

initial begin
    $display("Hello Verilog");
end

endmodule