`timescale 100ps / 100ps

module detector_010 (clk, reset, in, out);

// FILLME

endmodule
